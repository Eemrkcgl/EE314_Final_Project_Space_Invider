library verilog;
use verilog.vl_types.all;
entity enemy_vlg_vec_tst is
end enemy_vlg_vec_tst;
