library verilog;
use verilog.vl_types.all;
entity project_vlg_vec_tst is
end project_vlg_vec_tst;
